module plugin

fn test_plugin() {
	// stub
}
