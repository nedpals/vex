module vex

import server

pub fn server() server.Server{
	return server.server()
}