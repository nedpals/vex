module websocket

import x.websocket