module router

fn test_plugin() {
	// stub
}
